library verilog;
use verilog.vl_types.all;
entity roundKeyGen_vlg_vec_tst is
end roundKeyGen_vlg_vec_tst;
