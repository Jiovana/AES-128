library verilog;
use verilog.vl_types.all;
entity word_subBytes_vlg_vec_tst is
end word_subBytes_vlg_vec_tst;
